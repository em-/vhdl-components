package alu_operations is
    type ALU_OPERATION is (ADD, SUB, ADDS, SUBS, MULT, 
                        BITAND, BITOR, BITXOR,
                        FUNCLSL, FUNCLSR, FUNCRL, FUNCRR);
end alu_operations;
