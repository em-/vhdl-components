library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity multiplier is
    generic (N: integer := 4);
    port (A, B:     in  std_logic_vector (N-1 downto 0);
          O:        out std_logic_vector (2*N-1 downto 0)
    );
end multiplier;

architecture behavioral of multiplier is
begin
    O <= std_logic_vector(unsigned(unsigned(A) * unsigned(B)));
end behavioral;


architecture structural of multiplier is
    component fa
        port (A, B: in std_logic;
              Ci:   in  std_logic;
              S:    out std_logic;
              Co:   out std_logic);
    end component;
    component ha
        port (A, B:  in  std_logic;
              S, Co: out std_logic);
    end component;
    component and2
        port (A, B: in  std_logic;
              O:    out std_logic);
    end component;

    type SignalVector is array (N-1 downto 0) of std_logic_vector(N-1 downto 0);
    signal tAND, S, C: SignalVector;
begin
    ands: for i in B'Range generate
        ands_i: for j in A'Range generate
            ands_ij: and2 port map (B(i), A(j), tAND(i)(j));
        end generate;
    end generate;

    S(0) <= tAND(0);
    C(0) <= (others => '0');

    row: for i in 1 to N-1 generate
    O(i-1) <= S(i-1)(0);

    ha00: ha
    port map (S(i-1)(1), tAND(i)(0), S(i)(0), C(i)(0));
    fa01: fa
    port map (S(i-1)(2), tAND(i)(1), C(i)(0), S(i)(1), C(i)(1));
    fa02: fa
    port map (S(i-1)(3), tAND(i)(2), C(i)(1), S(i)(2), C(i)(2));
    fa03: fa
    port map (C(i-1)(3), tAND(i)(3), C(i)(2), S(i)(3), C(i)(3));
    end generate;

    O(6 downto 3) <= S(3);
    O(7) <= C(3)(3);
end structural;

configuration cfg_multiplier_behavioral of multiplier is
    for behavioral
    end for;
end cfg_multiplier_behavioral;

configuration cfg_multiplier_structural of multiplier is
    for structural
    end for;
end cfg_multiplier_structural;
